module bramki #(
    parameters
) (
    ports
);



endmodule